---
-- File: P3_PROG_START.vhd
-- Type: rtl_vhdl
-- Author: jellch
-- Created: 2025-11-28
-- Modified: 2025-11-28 02:22:25
-- Code_link: "[[rtl/boot/P3_PROG_START.vhd|P3_PROG_START.vhd]]"
-- Doc_link: "[[rtl/boot/P3_PROG_START.vhd.md|P3_PROG_START.vhd.md]]"
-- Self_link: "[[rtl/boot/P3_PROG_START.vhd|P3_PROG_START.vhd]]"
---


-- TODO: Add VHDL code here
-- This is a placeholder template for the .vhd file

-- See Also
-- ## [P3_PROG_START.vhd.md](rtl/boot/P3_PROG_START.vhd.md)
