---
-- File: L2_BUFF_LOADER.vhd
-- Type: rtl_vhdl
-- Author: jellch
-- Created: 2025-11-28
-- Modified: 2025-11-28 02:21:50
-- Code_link: "[[rtl/boot/L2_BUFF_LOADER.vhd|L2_BUFF_LOADER.vhd]]"
-- Doc_link: "[[rtl/boot/L2_BUFF_LOADER.vhd.md|L2_BUFF_LOADER.vhd.md]]"
-- Self_link: "[[rtl/boot/L2_BUFF_LOADER.vhd|L2_BUFF_LOADER.vhd]]"
---


-- TODO: Add VHDL code here
-- This is a placeholder template for the .vhd file

-- See Also
-- ## [L2_BUFF_LOADER.vhd.md](rtl/boot/L2_BUFF_LOADER.vhd.md)
