---
-- File: B0_BOOT_TOP.vhd
-- Type: rtl_vhdl
-- Author: jellch
-- Created: 2025-11-28
-- Modified: 2025-11-28 02:20:40
-- Code_link: "[[rtl/boot/B0_BOOT_TOP.vhd|B0_BOOT_TOP.vhd]]"
-- Doc_link: "[[rtl/boot/B0_BOOT_TOP.vhd.md|B0_BOOT_TOP.vhd.md]]"
-- Self_link: "[[rtl/boot/B0_BOOT_TOP.vhd|B0_BOOT_TOP.vhd]]"
---


-- TODO: Add VHDL code here
-- This is a placeholder template for the .vhd file

-- See Also
-- ## [B0_BOOT_TOP.vhd.md](rtl/boot/B0_BOOT_TOP.vhd.md)
